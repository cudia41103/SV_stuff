

package cache_types;
typedef enum logic [1:0] {
    way1 = 2'b00,
    way2 = 2'b01,
    way3 = 2'b10,
    way4 = 2'b11
}dmux_sel_t;
endpackage